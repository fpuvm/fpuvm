`ifndef AVALON_MM_MST_SEQUENCER
`define AVALON_MM_MST_SEQUENCER

class avalon_mm_mst_sequencer extends uvm_sequencer #(avalon_mm_xactn);
  `uvm_component_utils_begin (avalon_mm_mst_sequencer)
  `uvm_component_utils_end

  `FP_UVM_COMP_NEW
endclass : avalon_mm_mst_sequencer 

`endif //  AVALON_MM_MST_SEQUENCER


